magic
tech sky130A
magscale 1 2
timestamp 1670788656
<< obsli1 >>
rect 1104 2159 318872 437393
<< obsm1 >>
rect 106 2048 319410 437424
<< metal2 >>
rect 3974 439200 4030 440000
rect 6734 439200 6790 440000
rect 9494 439200 9550 440000
rect 12254 439200 12310 440000
rect 15014 439200 15070 440000
rect 17774 439200 17830 440000
rect 20534 439200 20590 440000
rect 23294 439200 23350 440000
rect 26054 439200 26110 440000
rect 28814 439200 28870 440000
rect 31574 439200 31630 440000
rect 34334 439200 34390 440000
rect 37094 439200 37150 440000
rect 39854 439200 39910 440000
rect 42614 439200 42670 440000
rect 45374 439200 45430 440000
rect 48134 439200 48190 440000
rect 50894 439200 50950 440000
rect 53654 439200 53710 440000
rect 56414 439200 56470 440000
rect 59174 439200 59230 440000
rect 61934 439200 61990 440000
rect 64694 439200 64750 440000
rect 67454 439200 67510 440000
rect 70214 439200 70270 440000
rect 72974 439200 73030 440000
rect 75734 439200 75790 440000
rect 78494 439200 78550 440000
rect 81254 439200 81310 440000
rect 84014 439200 84070 440000
rect 86774 439200 86830 440000
rect 89534 439200 89590 440000
rect 92294 439200 92350 440000
rect 95054 439200 95110 440000
rect 97814 439200 97870 440000
rect 100574 439200 100630 440000
rect 103334 439200 103390 440000
rect 106094 439200 106150 440000
rect 108854 439200 108910 440000
rect 111614 439200 111670 440000
rect 114374 439200 114430 440000
rect 117134 439200 117190 440000
rect 119894 439200 119950 440000
rect 122654 439200 122710 440000
rect 125414 439200 125470 440000
rect 128174 439200 128230 440000
rect 130934 439200 130990 440000
rect 133694 439200 133750 440000
rect 136454 439200 136510 440000
rect 139214 439200 139270 440000
rect 141974 439200 142030 440000
rect 144734 439200 144790 440000
rect 147494 439200 147550 440000
rect 150254 439200 150310 440000
rect 153014 439200 153070 440000
rect 155774 439200 155830 440000
rect 158534 439200 158590 440000
rect 161294 439200 161350 440000
rect 164054 439200 164110 440000
rect 166814 439200 166870 440000
rect 169574 439200 169630 440000
rect 172334 439200 172390 440000
rect 175094 439200 175150 440000
rect 177854 439200 177910 440000
rect 180614 439200 180670 440000
rect 183374 439200 183430 440000
rect 186134 439200 186190 440000
rect 188894 439200 188950 440000
rect 191654 439200 191710 440000
rect 194414 439200 194470 440000
rect 197174 439200 197230 440000
rect 199934 439200 199990 440000
rect 202694 439200 202750 440000
rect 205454 439200 205510 440000
rect 208214 439200 208270 440000
rect 210974 439200 211030 440000
rect 213734 439200 213790 440000
rect 216494 439200 216550 440000
rect 219254 439200 219310 440000
rect 222014 439200 222070 440000
rect 224774 439200 224830 440000
rect 227534 439200 227590 440000
rect 230294 439200 230350 440000
rect 233054 439200 233110 440000
rect 235814 439200 235870 440000
rect 238574 439200 238630 440000
rect 241334 439200 241390 440000
rect 244094 439200 244150 440000
rect 246854 439200 246910 440000
rect 249614 439200 249670 440000
rect 252374 439200 252430 440000
rect 255134 439200 255190 440000
rect 257894 439200 257950 440000
rect 260654 439200 260710 440000
rect 263414 439200 263470 440000
rect 266174 439200 266230 440000
rect 268934 439200 268990 440000
rect 271694 439200 271750 440000
rect 274454 439200 274510 440000
rect 277214 439200 277270 440000
rect 279974 439200 280030 440000
rect 282734 439200 282790 440000
rect 285494 439200 285550 440000
rect 288254 439200 288310 440000
rect 291014 439200 291070 440000
rect 293774 439200 293830 440000
rect 296534 439200 296590 440000
rect 299294 439200 299350 440000
rect 302054 439200 302110 440000
rect 304814 439200 304870 440000
rect 307574 439200 307630 440000
rect 310334 439200 310390 440000
rect 313094 439200 313150 440000
rect 315854 439200 315910 440000
rect 1490 0 1546 800
rect 2134 0 2190 800
rect 2778 0 2834 800
rect 3422 0 3478 800
rect 4066 0 4122 800
rect 4710 0 4766 800
rect 5354 0 5410 800
rect 5998 0 6054 800
rect 6642 0 6698 800
rect 7286 0 7342 800
rect 7930 0 7986 800
rect 8574 0 8630 800
rect 9218 0 9274 800
rect 9862 0 9918 800
rect 10506 0 10562 800
rect 11150 0 11206 800
rect 11794 0 11850 800
rect 12438 0 12494 800
rect 13082 0 13138 800
rect 13726 0 13782 800
rect 14370 0 14426 800
rect 15014 0 15070 800
rect 15658 0 15714 800
rect 16302 0 16358 800
rect 16946 0 17002 800
rect 17590 0 17646 800
rect 18234 0 18290 800
rect 18878 0 18934 800
rect 19522 0 19578 800
rect 20166 0 20222 800
rect 20810 0 20866 800
rect 21454 0 21510 800
rect 22098 0 22154 800
rect 22742 0 22798 800
rect 23386 0 23442 800
rect 24030 0 24086 800
rect 24674 0 24730 800
rect 25318 0 25374 800
rect 25962 0 26018 800
rect 26606 0 26662 800
rect 27250 0 27306 800
rect 27894 0 27950 800
rect 28538 0 28594 800
rect 29182 0 29238 800
rect 29826 0 29882 800
rect 30470 0 30526 800
rect 31114 0 31170 800
rect 31758 0 31814 800
rect 32402 0 32458 800
rect 33046 0 33102 800
rect 33690 0 33746 800
rect 34334 0 34390 800
rect 34978 0 35034 800
rect 35622 0 35678 800
rect 36266 0 36322 800
rect 36910 0 36966 800
rect 37554 0 37610 800
rect 38198 0 38254 800
rect 38842 0 38898 800
rect 39486 0 39542 800
rect 40130 0 40186 800
rect 40774 0 40830 800
rect 41418 0 41474 800
rect 42062 0 42118 800
rect 42706 0 42762 800
rect 43350 0 43406 800
rect 43994 0 44050 800
rect 44638 0 44694 800
rect 45282 0 45338 800
rect 45926 0 45982 800
rect 46570 0 46626 800
rect 47214 0 47270 800
rect 47858 0 47914 800
rect 48502 0 48558 800
rect 49146 0 49202 800
rect 49790 0 49846 800
rect 50434 0 50490 800
rect 51078 0 51134 800
rect 51722 0 51778 800
rect 52366 0 52422 800
rect 53010 0 53066 800
rect 53654 0 53710 800
rect 54298 0 54354 800
rect 54942 0 54998 800
rect 55586 0 55642 800
rect 56230 0 56286 800
rect 56874 0 56930 800
rect 57518 0 57574 800
rect 58162 0 58218 800
rect 58806 0 58862 800
rect 59450 0 59506 800
rect 60094 0 60150 800
rect 60738 0 60794 800
rect 61382 0 61438 800
rect 62026 0 62082 800
rect 62670 0 62726 800
rect 63314 0 63370 800
rect 63958 0 64014 800
rect 64602 0 64658 800
rect 65246 0 65302 800
rect 65890 0 65946 800
rect 66534 0 66590 800
rect 67178 0 67234 800
rect 67822 0 67878 800
rect 68466 0 68522 800
rect 69110 0 69166 800
rect 69754 0 69810 800
rect 70398 0 70454 800
rect 71042 0 71098 800
rect 71686 0 71742 800
rect 72330 0 72386 800
rect 72974 0 73030 800
rect 73618 0 73674 800
rect 74262 0 74318 800
rect 74906 0 74962 800
rect 75550 0 75606 800
rect 76194 0 76250 800
rect 76838 0 76894 800
rect 77482 0 77538 800
rect 78126 0 78182 800
rect 78770 0 78826 800
rect 79414 0 79470 800
rect 80058 0 80114 800
rect 80702 0 80758 800
rect 81346 0 81402 800
rect 81990 0 82046 800
rect 82634 0 82690 800
rect 83278 0 83334 800
rect 83922 0 83978 800
rect 84566 0 84622 800
rect 85210 0 85266 800
rect 85854 0 85910 800
rect 86498 0 86554 800
rect 87142 0 87198 800
rect 87786 0 87842 800
rect 88430 0 88486 800
rect 89074 0 89130 800
rect 89718 0 89774 800
rect 90362 0 90418 800
rect 91006 0 91062 800
rect 91650 0 91706 800
rect 92294 0 92350 800
rect 92938 0 92994 800
rect 93582 0 93638 800
rect 94226 0 94282 800
rect 94870 0 94926 800
rect 95514 0 95570 800
rect 96158 0 96214 800
rect 96802 0 96858 800
rect 97446 0 97502 800
rect 98090 0 98146 800
rect 98734 0 98790 800
rect 99378 0 99434 800
rect 100022 0 100078 800
rect 100666 0 100722 800
rect 101310 0 101366 800
rect 101954 0 102010 800
rect 102598 0 102654 800
rect 103242 0 103298 800
rect 103886 0 103942 800
rect 104530 0 104586 800
rect 105174 0 105230 800
rect 105818 0 105874 800
rect 106462 0 106518 800
rect 107106 0 107162 800
rect 107750 0 107806 800
rect 108394 0 108450 800
rect 109038 0 109094 800
rect 109682 0 109738 800
rect 110326 0 110382 800
rect 110970 0 111026 800
rect 111614 0 111670 800
rect 112258 0 112314 800
rect 112902 0 112958 800
rect 113546 0 113602 800
rect 114190 0 114246 800
rect 114834 0 114890 800
rect 115478 0 115534 800
rect 116122 0 116178 800
rect 116766 0 116822 800
rect 117410 0 117466 800
rect 118054 0 118110 800
rect 118698 0 118754 800
rect 119342 0 119398 800
rect 119986 0 120042 800
rect 120630 0 120686 800
rect 121274 0 121330 800
rect 121918 0 121974 800
rect 122562 0 122618 800
rect 123206 0 123262 800
rect 123850 0 123906 800
rect 124494 0 124550 800
rect 125138 0 125194 800
rect 125782 0 125838 800
rect 126426 0 126482 800
rect 127070 0 127126 800
rect 127714 0 127770 800
rect 128358 0 128414 800
rect 129002 0 129058 800
rect 129646 0 129702 800
rect 130290 0 130346 800
rect 130934 0 130990 800
rect 131578 0 131634 800
rect 132222 0 132278 800
rect 132866 0 132922 800
rect 133510 0 133566 800
rect 134154 0 134210 800
rect 134798 0 134854 800
rect 135442 0 135498 800
rect 136086 0 136142 800
rect 136730 0 136786 800
rect 137374 0 137430 800
rect 138018 0 138074 800
rect 138662 0 138718 800
rect 139306 0 139362 800
rect 139950 0 140006 800
rect 140594 0 140650 800
rect 141238 0 141294 800
rect 141882 0 141938 800
rect 142526 0 142582 800
rect 143170 0 143226 800
rect 143814 0 143870 800
rect 144458 0 144514 800
rect 145102 0 145158 800
rect 145746 0 145802 800
rect 146390 0 146446 800
rect 147034 0 147090 800
rect 147678 0 147734 800
rect 148322 0 148378 800
rect 148966 0 149022 800
rect 149610 0 149666 800
rect 150254 0 150310 800
rect 150898 0 150954 800
rect 151542 0 151598 800
rect 152186 0 152242 800
rect 152830 0 152886 800
rect 153474 0 153530 800
rect 154118 0 154174 800
rect 154762 0 154818 800
rect 155406 0 155462 800
rect 156050 0 156106 800
rect 156694 0 156750 800
rect 157338 0 157394 800
rect 157982 0 158038 800
rect 158626 0 158682 800
rect 159270 0 159326 800
rect 159914 0 159970 800
rect 160558 0 160614 800
rect 161202 0 161258 800
rect 161846 0 161902 800
rect 162490 0 162546 800
rect 163134 0 163190 800
rect 163778 0 163834 800
rect 164422 0 164478 800
rect 165066 0 165122 800
rect 165710 0 165766 800
rect 166354 0 166410 800
rect 166998 0 167054 800
rect 167642 0 167698 800
rect 168286 0 168342 800
rect 168930 0 168986 800
rect 169574 0 169630 800
rect 170218 0 170274 800
rect 170862 0 170918 800
rect 171506 0 171562 800
rect 172150 0 172206 800
rect 172794 0 172850 800
rect 173438 0 173494 800
rect 174082 0 174138 800
rect 174726 0 174782 800
rect 175370 0 175426 800
rect 176014 0 176070 800
rect 176658 0 176714 800
rect 177302 0 177358 800
rect 177946 0 178002 800
rect 178590 0 178646 800
rect 179234 0 179290 800
rect 179878 0 179934 800
rect 180522 0 180578 800
rect 181166 0 181222 800
rect 181810 0 181866 800
rect 182454 0 182510 800
rect 183098 0 183154 800
rect 183742 0 183798 800
rect 184386 0 184442 800
rect 185030 0 185086 800
rect 185674 0 185730 800
rect 186318 0 186374 800
rect 186962 0 187018 800
rect 187606 0 187662 800
rect 188250 0 188306 800
rect 188894 0 188950 800
rect 189538 0 189594 800
rect 190182 0 190238 800
rect 190826 0 190882 800
rect 191470 0 191526 800
rect 192114 0 192170 800
rect 192758 0 192814 800
rect 193402 0 193458 800
rect 194046 0 194102 800
rect 194690 0 194746 800
rect 195334 0 195390 800
rect 195978 0 196034 800
rect 196622 0 196678 800
rect 197266 0 197322 800
rect 197910 0 197966 800
rect 198554 0 198610 800
rect 199198 0 199254 800
rect 199842 0 199898 800
rect 200486 0 200542 800
rect 201130 0 201186 800
rect 201774 0 201830 800
rect 202418 0 202474 800
rect 203062 0 203118 800
rect 203706 0 203762 800
rect 204350 0 204406 800
rect 204994 0 205050 800
rect 205638 0 205694 800
rect 206282 0 206338 800
rect 206926 0 206982 800
rect 207570 0 207626 800
rect 208214 0 208270 800
rect 208858 0 208914 800
rect 209502 0 209558 800
rect 210146 0 210202 800
rect 210790 0 210846 800
rect 211434 0 211490 800
rect 212078 0 212134 800
rect 212722 0 212778 800
rect 213366 0 213422 800
rect 214010 0 214066 800
rect 214654 0 214710 800
rect 215298 0 215354 800
rect 215942 0 215998 800
rect 216586 0 216642 800
rect 217230 0 217286 800
rect 217874 0 217930 800
rect 218518 0 218574 800
rect 219162 0 219218 800
rect 219806 0 219862 800
rect 220450 0 220506 800
rect 221094 0 221150 800
rect 221738 0 221794 800
rect 222382 0 222438 800
rect 223026 0 223082 800
rect 223670 0 223726 800
rect 224314 0 224370 800
rect 224958 0 225014 800
rect 225602 0 225658 800
rect 226246 0 226302 800
rect 226890 0 226946 800
rect 227534 0 227590 800
rect 228178 0 228234 800
rect 228822 0 228878 800
rect 229466 0 229522 800
rect 230110 0 230166 800
rect 230754 0 230810 800
rect 231398 0 231454 800
rect 232042 0 232098 800
rect 232686 0 232742 800
rect 233330 0 233386 800
rect 233974 0 234030 800
rect 234618 0 234674 800
rect 235262 0 235318 800
rect 235906 0 235962 800
rect 236550 0 236606 800
rect 237194 0 237250 800
rect 237838 0 237894 800
rect 238482 0 238538 800
rect 239126 0 239182 800
rect 239770 0 239826 800
rect 240414 0 240470 800
rect 241058 0 241114 800
rect 241702 0 241758 800
rect 242346 0 242402 800
rect 242990 0 243046 800
rect 243634 0 243690 800
rect 244278 0 244334 800
rect 244922 0 244978 800
rect 245566 0 245622 800
rect 246210 0 246266 800
rect 246854 0 246910 800
rect 247498 0 247554 800
rect 248142 0 248198 800
rect 248786 0 248842 800
rect 249430 0 249486 800
rect 250074 0 250130 800
rect 250718 0 250774 800
rect 251362 0 251418 800
rect 252006 0 252062 800
rect 252650 0 252706 800
rect 253294 0 253350 800
rect 253938 0 253994 800
rect 254582 0 254638 800
rect 255226 0 255282 800
rect 255870 0 255926 800
rect 256514 0 256570 800
rect 257158 0 257214 800
rect 257802 0 257858 800
rect 258446 0 258502 800
rect 259090 0 259146 800
rect 259734 0 259790 800
rect 260378 0 260434 800
rect 261022 0 261078 800
rect 261666 0 261722 800
rect 262310 0 262366 800
rect 262954 0 263010 800
rect 263598 0 263654 800
rect 264242 0 264298 800
rect 264886 0 264942 800
rect 265530 0 265586 800
rect 266174 0 266230 800
rect 266818 0 266874 800
rect 267462 0 267518 800
rect 268106 0 268162 800
rect 268750 0 268806 800
rect 269394 0 269450 800
rect 270038 0 270094 800
rect 270682 0 270738 800
rect 271326 0 271382 800
rect 271970 0 272026 800
rect 272614 0 272670 800
rect 273258 0 273314 800
rect 273902 0 273958 800
rect 274546 0 274602 800
rect 275190 0 275246 800
rect 275834 0 275890 800
rect 276478 0 276534 800
rect 277122 0 277178 800
rect 277766 0 277822 800
rect 278410 0 278466 800
rect 279054 0 279110 800
rect 279698 0 279754 800
rect 280342 0 280398 800
rect 280986 0 281042 800
rect 281630 0 281686 800
rect 282274 0 282330 800
rect 282918 0 282974 800
rect 283562 0 283618 800
rect 284206 0 284262 800
rect 284850 0 284906 800
rect 285494 0 285550 800
rect 286138 0 286194 800
rect 286782 0 286838 800
rect 287426 0 287482 800
rect 288070 0 288126 800
rect 288714 0 288770 800
rect 289358 0 289414 800
rect 290002 0 290058 800
rect 290646 0 290702 800
rect 291290 0 291346 800
rect 291934 0 291990 800
rect 292578 0 292634 800
rect 293222 0 293278 800
rect 293866 0 293922 800
rect 294510 0 294566 800
rect 295154 0 295210 800
rect 295798 0 295854 800
rect 296442 0 296498 800
rect 297086 0 297142 800
rect 297730 0 297786 800
rect 298374 0 298430 800
rect 299018 0 299074 800
rect 299662 0 299718 800
rect 300306 0 300362 800
rect 300950 0 301006 800
rect 301594 0 301650 800
rect 302238 0 302294 800
rect 302882 0 302938 800
rect 303526 0 303582 800
rect 304170 0 304226 800
rect 304814 0 304870 800
rect 305458 0 305514 800
rect 306102 0 306158 800
rect 306746 0 306802 800
rect 307390 0 307446 800
rect 308034 0 308090 800
rect 308678 0 308734 800
rect 309322 0 309378 800
rect 309966 0 310022 800
rect 310610 0 310666 800
rect 311254 0 311310 800
rect 311898 0 311954 800
rect 312542 0 312598 800
rect 313186 0 313242 800
rect 313830 0 313886 800
rect 314474 0 314530 800
rect 315118 0 315174 800
rect 315762 0 315818 800
rect 316406 0 316462 800
rect 317050 0 317106 800
rect 317694 0 317750 800
rect 318338 0 318394 800
<< obsm2 >>
rect 112 439144 3918 439362
rect 4086 439144 6678 439362
rect 6846 439144 9438 439362
rect 9606 439144 12198 439362
rect 12366 439144 14958 439362
rect 15126 439144 17718 439362
rect 17886 439144 20478 439362
rect 20646 439144 23238 439362
rect 23406 439144 25998 439362
rect 26166 439144 28758 439362
rect 28926 439144 31518 439362
rect 31686 439144 34278 439362
rect 34446 439144 37038 439362
rect 37206 439144 39798 439362
rect 39966 439144 42558 439362
rect 42726 439144 45318 439362
rect 45486 439144 48078 439362
rect 48246 439144 50838 439362
rect 51006 439144 53598 439362
rect 53766 439144 56358 439362
rect 56526 439144 59118 439362
rect 59286 439144 61878 439362
rect 62046 439144 64638 439362
rect 64806 439144 67398 439362
rect 67566 439144 70158 439362
rect 70326 439144 72918 439362
rect 73086 439144 75678 439362
rect 75846 439144 78438 439362
rect 78606 439144 81198 439362
rect 81366 439144 83958 439362
rect 84126 439144 86718 439362
rect 86886 439144 89478 439362
rect 89646 439144 92238 439362
rect 92406 439144 94998 439362
rect 95166 439144 97758 439362
rect 97926 439144 100518 439362
rect 100686 439144 103278 439362
rect 103446 439144 106038 439362
rect 106206 439144 108798 439362
rect 108966 439144 111558 439362
rect 111726 439144 114318 439362
rect 114486 439144 117078 439362
rect 117246 439144 119838 439362
rect 120006 439144 122598 439362
rect 122766 439144 125358 439362
rect 125526 439144 128118 439362
rect 128286 439144 130878 439362
rect 131046 439144 133638 439362
rect 133806 439144 136398 439362
rect 136566 439144 139158 439362
rect 139326 439144 141918 439362
rect 142086 439144 144678 439362
rect 144846 439144 147438 439362
rect 147606 439144 150198 439362
rect 150366 439144 152958 439362
rect 153126 439144 155718 439362
rect 155886 439144 158478 439362
rect 158646 439144 161238 439362
rect 161406 439144 163998 439362
rect 164166 439144 166758 439362
rect 166926 439144 169518 439362
rect 169686 439144 172278 439362
rect 172446 439144 175038 439362
rect 175206 439144 177798 439362
rect 177966 439144 180558 439362
rect 180726 439144 183318 439362
rect 183486 439144 186078 439362
rect 186246 439144 188838 439362
rect 189006 439144 191598 439362
rect 191766 439144 194358 439362
rect 194526 439144 197118 439362
rect 197286 439144 199878 439362
rect 200046 439144 202638 439362
rect 202806 439144 205398 439362
rect 205566 439144 208158 439362
rect 208326 439144 210918 439362
rect 211086 439144 213678 439362
rect 213846 439144 216438 439362
rect 216606 439144 219198 439362
rect 219366 439144 221958 439362
rect 222126 439144 224718 439362
rect 224886 439144 227478 439362
rect 227646 439144 230238 439362
rect 230406 439144 232998 439362
rect 233166 439144 235758 439362
rect 235926 439144 238518 439362
rect 238686 439144 241278 439362
rect 241446 439144 244038 439362
rect 244206 439144 246798 439362
rect 246966 439144 249558 439362
rect 249726 439144 252318 439362
rect 252486 439144 255078 439362
rect 255246 439144 257838 439362
rect 258006 439144 260598 439362
rect 260766 439144 263358 439362
rect 263526 439144 266118 439362
rect 266286 439144 268878 439362
rect 269046 439144 271638 439362
rect 271806 439144 274398 439362
rect 274566 439144 277158 439362
rect 277326 439144 279918 439362
rect 280086 439144 282678 439362
rect 282846 439144 285438 439362
rect 285606 439144 288198 439362
rect 288366 439144 290958 439362
rect 291126 439144 293718 439362
rect 293886 439144 296478 439362
rect 296646 439144 299238 439362
rect 299406 439144 301998 439362
rect 302166 439144 304758 439362
rect 304926 439144 307518 439362
rect 307686 439144 310278 439362
rect 310446 439144 313038 439362
rect 313206 439144 315798 439362
rect 315966 439144 319404 439362
rect 112 856 319404 439144
rect 112 800 1434 856
rect 1602 800 2078 856
rect 2246 800 2722 856
rect 2890 800 3366 856
rect 3534 800 4010 856
rect 4178 800 4654 856
rect 4822 800 5298 856
rect 5466 800 5942 856
rect 6110 800 6586 856
rect 6754 800 7230 856
rect 7398 800 7874 856
rect 8042 800 8518 856
rect 8686 800 9162 856
rect 9330 800 9806 856
rect 9974 800 10450 856
rect 10618 800 11094 856
rect 11262 800 11738 856
rect 11906 800 12382 856
rect 12550 800 13026 856
rect 13194 800 13670 856
rect 13838 800 14314 856
rect 14482 800 14958 856
rect 15126 800 15602 856
rect 15770 800 16246 856
rect 16414 800 16890 856
rect 17058 800 17534 856
rect 17702 800 18178 856
rect 18346 800 18822 856
rect 18990 800 19466 856
rect 19634 800 20110 856
rect 20278 800 20754 856
rect 20922 800 21398 856
rect 21566 800 22042 856
rect 22210 800 22686 856
rect 22854 800 23330 856
rect 23498 800 23974 856
rect 24142 800 24618 856
rect 24786 800 25262 856
rect 25430 800 25906 856
rect 26074 800 26550 856
rect 26718 800 27194 856
rect 27362 800 27838 856
rect 28006 800 28482 856
rect 28650 800 29126 856
rect 29294 800 29770 856
rect 29938 800 30414 856
rect 30582 800 31058 856
rect 31226 800 31702 856
rect 31870 800 32346 856
rect 32514 800 32990 856
rect 33158 800 33634 856
rect 33802 800 34278 856
rect 34446 800 34922 856
rect 35090 800 35566 856
rect 35734 800 36210 856
rect 36378 800 36854 856
rect 37022 800 37498 856
rect 37666 800 38142 856
rect 38310 800 38786 856
rect 38954 800 39430 856
rect 39598 800 40074 856
rect 40242 800 40718 856
rect 40886 800 41362 856
rect 41530 800 42006 856
rect 42174 800 42650 856
rect 42818 800 43294 856
rect 43462 800 43938 856
rect 44106 800 44582 856
rect 44750 800 45226 856
rect 45394 800 45870 856
rect 46038 800 46514 856
rect 46682 800 47158 856
rect 47326 800 47802 856
rect 47970 800 48446 856
rect 48614 800 49090 856
rect 49258 800 49734 856
rect 49902 800 50378 856
rect 50546 800 51022 856
rect 51190 800 51666 856
rect 51834 800 52310 856
rect 52478 800 52954 856
rect 53122 800 53598 856
rect 53766 800 54242 856
rect 54410 800 54886 856
rect 55054 800 55530 856
rect 55698 800 56174 856
rect 56342 800 56818 856
rect 56986 800 57462 856
rect 57630 800 58106 856
rect 58274 800 58750 856
rect 58918 800 59394 856
rect 59562 800 60038 856
rect 60206 800 60682 856
rect 60850 800 61326 856
rect 61494 800 61970 856
rect 62138 800 62614 856
rect 62782 800 63258 856
rect 63426 800 63902 856
rect 64070 800 64546 856
rect 64714 800 65190 856
rect 65358 800 65834 856
rect 66002 800 66478 856
rect 66646 800 67122 856
rect 67290 800 67766 856
rect 67934 800 68410 856
rect 68578 800 69054 856
rect 69222 800 69698 856
rect 69866 800 70342 856
rect 70510 800 70986 856
rect 71154 800 71630 856
rect 71798 800 72274 856
rect 72442 800 72918 856
rect 73086 800 73562 856
rect 73730 800 74206 856
rect 74374 800 74850 856
rect 75018 800 75494 856
rect 75662 800 76138 856
rect 76306 800 76782 856
rect 76950 800 77426 856
rect 77594 800 78070 856
rect 78238 800 78714 856
rect 78882 800 79358 856
rect 79526 800 80002 856
rect 80170 800 80646 856
rect 80814 800 81290 856
rect 81458 800 81934 856
rect 82102 800 82578 856
rect 82746 800 83222 856
rect 83390 800 83866 856
rect 84034 800 84510 856
rect 84678 800 85154 856
rect 85322 800 85798 856
rect 85966 800 86442 856
rect 86610 800 87086 856
rect 87254 800 87730 856
rect 87898 800 88374 856
rect 88542 800 89018 856
rect 89186 800 89662 856
rect 89830 800 90306 856
rect 90474 800 90950 856
rect 91118 800 91594 856
rect 91762 800 92238 856
rect 92406 800 92882 856
rect 93050 800 93526 856
rect 93694 800 94170 856
rect 94338 800 94814 856
rect 94982 800 95458 856
rect 95626 800 96102 856
rect 96270 800 96746 856
rect 96914 800 97390 856
rect 97558 800 98034 856
rect 98202 800 98678 856
rect 98846 800 99322 856
rect 99490 800 99966 856
rect 100134 800 100610 856
rect 100778 800 101254 856
rect 101422 800 101898 856
rect 102066 800 102542 856
rect 102710 800 103186 856
rect 103354 800 103830 856
rect 103998 800 104474 856
rect 104642 800 105118 856
rect 105286 800 105762 856
rect 105930 800 106406 856
rect 106574 800 107050 856
rect 107218 800 107694 856
rect 107862 800 108338 856
rect 108506 800 108982 856
rect 109150 800 109626 856
rect 109794 800 110270 856
rect 110438 800 110914 856
rect 111082 800 111558 856
rect 111726 800 112202 856
rect 112370 800 112846 856
rect 113014 800 113490 856
rect 113658 800 114134 856
rect 114302 800 114778 856
rect 114946 800 115422 856
rect 115590 800 116066 856
rect 116234 800 116710 856
rect 116878 800 117354 856
rect 117522 800 117998 856
rect 118166 800 118642 856
rect 118810 800 119286 856
rect 119454 800 119930 856
rect 120098 800 120574 856
rect 120742 800 121218 856
rect 121386 800 121862 856
rect 122030 800 122506 856
rect 122674 800 123150 856
rect 123318 800 123794 856
rect 123962 800 124438 856
rect 124606 800 125082 856
rect 125250 800 125726 856
rect 125894 800 126370 856
rect 126538 800 127014 856
rect 127182 800 127658 856
rect 127826 800 128302 856
rect 128470 800 128946 856
rect 129114 800 129590 856
rect 129758 800 130234 856
rect 130402 800 130878 856
rect 131046 800 131522 856
rect 131690 800 132166 856
rect 132334 800 132810 856
rect 132978 800 133454 856
rect 133622 800 134098 856
rect 134266 800 134742 856
rect 134910 800 135386 856
rect 135554 800 136030 856
rect 136198 800 136674 856
rect 136842 800 137318 856
rect 137486 800 137962 856
rect 138130 800 138606 856
rect 138774 800 139250 856
rect 139418 800 139894 856
rect 140062 800 140538 856
rect 140706 800 141182 856
rect 141350 800 141826 856
rect 141994 800 142470 856
rect 142638 800 143114 856
rect 143282 800 143758 856
rect 143926 800 144402 856
rect 144570 800 145046 856
rect 145214 800 145690 856
rect 145858 800 146334 856
rect 146502 800 146978 856
rect 147146 800 147622 856
rect 147790 800 148266 856
rect 148434 800 148910 856
rect 149078 800 149554 856
rect 149722 800 150198 856
rect 150366 800 150842 856
rect 151010 800 151486 856
rect 151654 800 152130 856
rect 152298 800 152774 856
rect 152942 800 153418 856
rect 153586 800 154062 856
rect 154230 800 154706 856
rect 154874 800 155350 856
rect 155518 800 155994 856
rect 156162 800 156638 856
rect 156806 800 157282 856
rect 157450 800 157926 856
rect 158094 800 158570 856
rect 158738 800 159214 856
rect 159382 800 159858 856
rect 160026 800 160502 856
rect 160670 800 161146 856
rect 161314 800 161790 856
rect 161958 800 162434 856
rect 162602 800 163078 856
rect 163246 800 163722 856
rect 163890 800 164366 856
rect 164534 800 165010 856
rect 165178 800 165654 856
rect 165822 800 166298 856
rect 166466 800 166942 856
rect 167110 800 167586 856
rect 167754 800 168230 856
rect 168398 800 168874 856
rect 169042 800 169518 856
rect 169686 800 170162 856
rect 170330 800 170806 856
rect 170974 800 171450 856
rect 171618 800 172094 856
rect 172262 800 172738 856
rect 172906 800 173382 856
rect 173550 800 174026 856
rect 174194 800 174670 856
rect 174838 800 175314 856
rect 175482 800 175958 856
rect 176126 800 176602 856
rect 176770 800 177246 856
rect 177414 800 177890 856
rect 178058 800 178534 856
rect 178702 800 179178 856
rect 179346 800 179822 856
rect 179990 800 180466 856
rect 180634 800 181110 856
rect 181278 800 181754 856
rect 181922 800 182398 856
rect 182566 800 183042 856
rect 183210 800 183686 856
rect 183854 800 184330 856
rect 184498 800 184974 856
rect 185142 800 185618 856
rect 185786 800 186262 856
rect 186430 800 186906 856
rect 187074 800 187550 856
rect 187718 800 188194 856
rect 188362 800 188838 856
rect 189006 800 189482 856
rect 189650 800 190126 856
rect 190294 800 190770 856
rect 190938 800 191414 856
rect 191582 800 192058 856
rect 192226 800 192702 856
rect 192870 800 193346 856
rect 193514 800 193990 856
rect 194158 800 194634 856
rect 194802 800 195278 856
rect 195446 800 195922 856
rect 196090 800 196566 856
rect 196734 800 197210 856
rect 197378 800 197854 856
rect 198022 800 198498 856
rect 198666 800 199142 856
rect 199310 800 199786 856
rect 199954 800 200430 856
rect 200598 800 201074 856
rect 201242 800 201718 856
rect 201886 800 202362 856
rect 202530 800 203006 856
rect 203174 800 203650 856
rect 203818 800 204294 856
rect 204462 800 204938 856
rect 205106 800 205582 856
rect 205750 800 206226 856
rect 206394 800 206870 856
rect 207038 800 207514 856
rect 207682 800 208158 856
rect 208326 800 208802 856
rect 208970 800 209446 856
rect 209614 800 210090 856
rect 210258 800 210734 856
rect 210902 800 211378 856
rect 211546 800 212022 856
rect 212190 800 212666 856
rect 212834 800 213310 856
rect 213478 800 213954 856
rect 214122 800 214598 856
rect 214766 800 215242 856
rect 215410 800 215886 856
rect 216054 800 216530 856
rect 216698 800 217174 856
rect 217342 800 217818 856
rect 217986 800 218462 856
rect 218630 800 219106 856
rect 219274 800 219750 856
rect 219918 800 220394 856
rect 220562 800 221038 856
rect 221206 800 221682 856
rect 221850 800 222326 856
rect 222494 800 222970 856
rect 223138 800 223614 856
rect 223782 800 224258 856
rect 224426 800 224902 856
rect 225070 800 225546 856
rect 225714 800 226190 856
rect 226358 800 226834 856
rect 227002 800 227478 856
rect 227646 800 228122 856
rect 228290 800 228766 856
rect 228934 800 229410 856
rect 229578 800 230054 856
rect 230222 800 230698 856
rect 230866 800 231342 856
rect 231510 800 231986 856
rect 232154 800 232630 856
rect 232798 800 233274 856
rect 233442 800 233918 856
rect 234086 800 234562 856
rect 234730 800 235206 856
rect 235374 800 235850 856
rect 236018 800 236494 856
rect 236662 800 237138 856
rect 237306 800 237782 856
rect 237950 800 238426 856
rect 238594 800 239070 856
rect 239238 800 239714 856
rect 239882 800 240358 856
rect 240526 800 241002 856
rect 241170 800 241646 856
rect 241814 800 242290 856
rect 242458 800 242934 856
rect 243102 800 243578 856
rect 243746 800 244222 856
rect 244390 800 244866 856
rect 245034 800 245510 856
rect 245678 800 246154 856
rect 246322 800 246798 856
rect 246966 800 247442 856
rect 247610 800 248086 856
rect 248254 800 248730 856
rect 248898 800 249374 856
rect 249542 800 250018 856
rect 250186 800 250662 856
rect 250830 800 251306 856
rect 251474 800 251950 856
rect 252118 800 252594 856
rect 252762 800 253238 856
rect 253406 800 253882 856
rect 254050 800 254526 856
rect 254694 800 255170 856
rect 255338 800 255814 856
rect 255982 800 256458 856
rect 256626 800 257102 856
rect 257270 800 257746 856
rect 257914 800 258390 856
rect 258558 800 259034 856
rect 259202 800 259678 856
rect 259846 800 260322 856
rect 260490 800 260966 856
rect 261134 800 261610 856
rect 261778 800 262254 856
rect 262422 800 262898 856
rect 263066 800 263542 856
rect 263710 800 264186 856
rect 264354 800 264830 856
rect 264998 800 265474 856
rect 265642 800 266118 856
rect 266286 800 266762 856
rect 266930 800 267406 856
rect 267574 800 268050 856
rect 268218 800 268694 856
rect 268862 800 269338 856
rect 269506 800 269982 856
rect 270150 800 270626 856
rect 270794 800 271270 856
rect 271438 800 271914 856
rect 272082 800 272558 856
rect 272726 800 273202 856
rect 273370 800 273846 856
rect 274014 800 274490 856
rect 274658 800 275134 856
rect 275302 800 275778 856
rect 275946 800 276422 856
rect 276590 800 277066 856
rect 277234 800 277710 856
rect 277878 800 278354 856
rect 278522 800 278998 856
rect 279166 800 279642 856
rect 279810 800 280286 856
rect 280454 800 280930 856
rect 281098 800 281574 856
rect 281742 800 282218 856
rect 282386 800 282862 856
rect 283030 800 283506 856
rect 283674 800 284150 856
rect 284318 800 284794 856
rect 284962 800 285438 856
rect 285606 800 286082 856
rect 286250 800 286726 856
rect 286894 800 287370 856
rect 287538 800 288014 856
rect 288182 800 288658 856
rect 288826 800 289302 856
rect 289470 800 289946 856
rect 290114 800 290590 856
rect 290758 800 291234 856
rect 291402 800 291878 856
rect 292046 800 292522 856
rect 292690 800 293166 856
rect 293334 800 293810 856
rect 293978 800 294454 856
rect 294622 800 295098 856
rect 295266 800 295742 856
rect 295910 800 296386 856
rect 296554 800 297030 856
rect 297198 800 297674 856
rect 297842 800 298318 856
rect 298486 800 298962 856
rect 299130 800 299606 856
rect 299774 800 300250 856
rect 300418 800 300894 856
rect 301062 800 301538 856
rect 301706 800 302182 856
rect 302350 800 302826 856
rect 302994 800 303470 856
rect 303638 800 304114 856
rect 304282 800 304758 856
rect 304926 800 305402 856
rect 305570 800 306046 856
rect 306214 800 306690 856
rect 306858 800 307334 856
rect 307502 800 307978 856
rect 308146 800 308622 856
rect 308790 800 309266 856
rect 309434 800 309910 856
rect 310078 800 310554 856
rect 310722 800 311198 856
rect 311366 800 311842 856
rect 312010 800 312486 856
rect 312654 800 313130 856
rect 313298 800 313774 856
rect 313942 800 314418 856
rect 314586 800 315062 856
rect 315230 800 315706 856
rect 315874 800 316350 856
rect 316518 800 316994 856
rect 317162 800 317638 856
rect 317806 800 318282 856
rect 318450 800 319404 856
<< obsm3 >>
rect 197 2143 319227 437409
<< metal4 >>
rect 4208 2128 4528 437424
rect 19568 2128 19888 437424
rect 34928 2128 35248 437424
rect 50288 2128 50608 437424
rect 65648 2128 65968 437424
rect 81008 2128 81328 437424
rect 96368 2128 96688 437424
rect 111728 2128 112048 437424
rect 127088 2128 127408 437424
rect 142448 2128 142768 437424
rect 157808 2128 158128 437424
rect 173168 2128 173488 437424
rect 188528 2128 188848 437424
rect 203888 2128 204208 437424
rect 219248 2128 219568 437424
rect 234608 2128 234928 437424
rect 249968 2128 250288 437424
rect 265328 2128 265648 437424
rect 280688 2128 281008 437424
rect 296048 2128 296368 437424
rect 311408 2128 311728 437424
<< obsm4 >>
rect 243 2347 4128 437069
rect 4608 2347 19488 437069
rect 19968 2347 34848 437069
rect 35328 2347 50208 437069
rect 50688 2347 65568 437069
rect 66048 2347 80928 437069
rect 81408 2347 96288 437069
rect 96768 2347 111648 437069
rect 112128 2347 127008 437069
rect 127488 2347 142368 437069
rect 142848 2347 157728 437069
rect 158208 2347 173088 437069
rect 173568 2347 188448 437069
rect 188928 2347 203808 437069
rect 204288 2347 219168 437069
rect 219648 2347 234528 437069
rect 235008 2347 249888 437069
rect 250368 2347 265248 437069
rect 265728 2347 280608 437069
rect 281088 2347 295968 437069
rect 296448 2347 311328 437069
rect 311808 2347 316605 437069
<< labels >>
rlabel metal2 s 3974 439200 4030 440000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 86774 439200 86830 440000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 95054 439200 95110 440000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 103334 439200 103390 440000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 111614 439200 111670 440000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 119894 439200 119950 440000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 128174 439200 128230 440000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 136454 439200 136510 440000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 144734 439200 144790 440000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 153014 439200 153070 440000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 161294 439200 161350 440000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 12254 439200 12310 440000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 169574 439200 169630 440000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 177854 439200 177910 440000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 186134 439200 186190 440000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 194414 439200 194470 440000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 202694 439200 202750 440000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 210974 439200 211030 440000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 219254 439200 219310 440000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 227534 439200 227590 440000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 235814 439200 235870 440000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 244094 439200 244150 440000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 20534 439200 20590 440000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 252374 439200 252430 440000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 260654 439200 260710 440000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 268934 439200 268990 440000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 277214 439200 277270 440000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 285494 439200 285550 440000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 293774 439200 293830 440000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 302054 439200 302110 440000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 310334 439200 310390 440000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 28814 439200 28870 440000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 37094 439200 37150 440000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 45374 439200 45430 440000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 53654 439200 53710 440000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 61934 439200 61990 440000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 70214 439200 70270 440000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 78494 439200 78550 440000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 6734 439200 6790 440000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 89534 439200 89590 440000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 97814 439200 97870 440000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 106094 439200 106150 440000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 114374 439200 114430 440000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 122654 439200 122710 440000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 130934 439200 130990 440000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 139214 439200 139270 440000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 147494 439200 147550 440000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 155774 439200 155830 440000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 164054 439200 164110 440000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 15014 439200 15070 440000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 172334 439200 172390 440000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 180614 439200 180670 440000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 188894 439200 188950 440000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 197174 439200 197230 440000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 205454 439200 205510 440000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 213734 439200 213790 440000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 222014 439200 222070 440000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 230294 439200 230350 440000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 238574 439200 238630 440000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 246854 439200 246910 440000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 23294 439200 23350 440000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 255134 439200 255190 440000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 263414 439200 263470 440000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 271694 439200 271750 440000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 279974 439200 280030 440000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 288254 439200 288310 440000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 296534 439200 296590 440000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 304814 439200 304870 440000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 313094 439200 313150 440000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 31574 439200 31630 440000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 39854 439200 39910 440000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 48134 439200 48190 440000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 56414 439200 56470 440000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 64694 439200 64750 440000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 72974 439200 73030 440000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 81254 439200 81310 440000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 9494 439200 9550 440000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 92294 439200 92350 440000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 100574 439200 100630 440000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 108854 439200 108910 440000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 117134 439200 117190 440000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 125414 439200 125470 440000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 133694 439200 133750 440000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 141974 439200 142030 440000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 150254 439200 150310 440000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 158534 439200 158590 440000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 166814 439200 166870 440000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 17774 439200 17830 440000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 175094 439200 175150 440000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 183374 439200 183430 440000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 191654 439200 191710 440000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 199934 439200 199990 440000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 208214 439200 208270 440000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 216494 439200 216550 440000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 224774 439200 224830 440000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 233054 439200 233110 440000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 241334 439200 241390 440000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 249614 439200 249670 440000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 26054 439200 26110 440000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 257894 439200 257950 440000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 266174 439200 266230 440000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 274454 439200 274510 440000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 282734 439200 282790 440000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 291014 439200 291070 440000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 299294 439200 299350 440000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 307574 439200 307630 440000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 315854 439200 315910 440000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 34334 439200 34390 440000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 42614 439200 42670 440000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 50894 439200 50950 440000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 59174 439200 59230 440000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 67454 439200 67510 440000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 75734 439200 75790 440000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 84014 439200 84070 440000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 317050 0 317106 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 317694 0 317750 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 318338 0 318394 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 262954 0 263010 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 264886 0 264942 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 266818 0 266874 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 268750 0 268806 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 270682 0 270738 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 272614 0 272670 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 274546 0 274602 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 276478 0 276534 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 278410 0 278466 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 280342 0 280398 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 282274 0 282330 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 284206 0 284262 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 286138 0 286194 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 288070 0 288126 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 290002 0 290058 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 291934 0 291990 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 293866 0 293922 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 295798 0 295854 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 297730 0 297786 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 299662 0 299718 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 301594 0 301650 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 303526 0 303582 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 305458 0 305514 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 307390 0 307446 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 309322 0 309378 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 311254 0 311310 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 313186 0 313242 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 315118 0 315174 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 176014 0 176070 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 179878 0 179934 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 181810 0 181866 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 185674 0 185730 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 187606 0 187662 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 191470 0 191526 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 193402 0 193458 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 195334 0 195390 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 197266 0 197322 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 199198 0 199254 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 201130 0 201186 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 204994 0 205050 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 206926 0 206982 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 208858 0 208914 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 210790 0 210846 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 212722 0 212778 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 214654 0 214710 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 216586 0 216642 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 218518 0 218574 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 220450 0 220506 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 222382 0 222438 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 224314 0 224370 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 226246 0 226302 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 228178 0 228234 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 230110 0 230166 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 232042 0 232098 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 233974 0 234030 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 235906 0 235962 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 237838 0 237894 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 239770 0 239826 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 243634 0 243690 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 247498 0 247554 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 249430 0 249486 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 251362 0 251418 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 253294 0 253350 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 255226 0 255282 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 257158 0 257214 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 259090 0 259146 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 261022 0 261078 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 263598 0 263654 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 265530 0 265586 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 267462 0 267518 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 269394 0 269450 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 271326 0 271382 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 273258 0 273314 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 275190 0 275246 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 277122 0 277178 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 279054 0 279110 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 280986 0 281042 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 282918 0 282974 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 284850 0 284906 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 286782 0 286838 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 288714 0 288770 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 290646 0 290702 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 292578 0 292634 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 294510 0 294566 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 296442 0 296498 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 298374 0 298430 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 300306 0 300362 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 302238 0 302294 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 304170 0 304226 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 306102 0 306158 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 308034 0 308090 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 309966 0 310022 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 311898 0 311954 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 313830 0 313886 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 315762 0 315818 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 95514 0 95570 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 97446 0 97502 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 103242 0 103298 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 105174 0 105230 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 120630 0 120686 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 122562 0 122618 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 128358 0 128414 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 132222 0 132278 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 145746 0 145802 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 147678 0 147734 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 151542 0 151598 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 153474 0 153530 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 159270 0 159326 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 163134 0 163190 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 165066 0 165122 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 166998 0 167054 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 170862 0 170918 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 172794 0 172850 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 174726 0 174782 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 176658 0 176714 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 178590 0 178646 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 180522 0 180578 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 182454 0 182510 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 184386 0 184442 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 186318 0 186374 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 188250 0 188306 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 190182 0 190238 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 192114 0 192170 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 194046 0 194102 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 195978 0 196034 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 197910 0 197966 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 199842 0 199898 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 201774 0 201830 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 203706 0 203762 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 205638 0 205694 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 207570 0 207626 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 209502 0 209558 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 211434 0 211490 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 213366 0 213422 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 215298 0 215354 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 217230 0 217286 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 219162 0 219218 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 221094 0 221150 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 223026 0 223082 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 224958 0 225014 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 226890 0 226946 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 228822 0 228878 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 230754 0 230810 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 232686 0 232742 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 234618 0 234674 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 236550 0 236606 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 238482 0 238538 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 240414 0 240470 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 242346 0 242402 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 244278 0 244334 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 246210 0 246266 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 248142 0 248198 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 250074 0 250130 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 252006 0 252062 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 253938 0 253994 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 255870 0 255926 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 257802 0 257858 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 259734 0 259790 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 261666 0 261722 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 264242 0 264298 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 266174 0 266230 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 268106 0 268162 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 270038 0 270094 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 271970 0 272026 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 273902 0 273958 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 275834 0 275890 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 277766 0 277822 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 279698 0 279754 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 281630 0 281686 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 283562 0 283618 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 285494 0 285550 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 287426 0 287482 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 289358 0 289414 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 291290 0 291346 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 293222 0 293278 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 295154 0 295210 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 297086 0 297142 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 299018 0 299074 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 300950 0 301006 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 302882 0 302938 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 304814 0 304870 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 306746 0 306802 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 308678 0 308734 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 310610 0 310666 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 312542 0 312598 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 314474 0 314530 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 316406 0 316462 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 132866 0 132922 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 169574 0 169630 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 173438 0 173494 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 179234 0 179290 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 181166 0 181222 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 185030 0 185086 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 188894 0 188950 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 192758 0 192814 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 194690 0 194746 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 196622 0 196678 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 200486 0 200542 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 202418 0 202474 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 204350 0 204406 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 206282 0 206338 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 208214 0 208270 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 210146 0 210202 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 212078 0 212134 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 214010 0 214066 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 215942 0 215998 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 217874 0 217930 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 219806 0 219862 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 221738 0 221794 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 223670 0 223726 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 225602 0 225658 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 227534 0 227590 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 229466 0 229522 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 231398 0 231454 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 233330 0 233386 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 235262 0 235318 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 237194 0 237250 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 239126 0 239182 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 241058 0 241114 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 242990 0 243046 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 244922 0 244978 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 246854 0 246910 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 248786 0 248842 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 250718 0 250774 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 252650 0 252706 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 254582 0 254638 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 256514 0 256570 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 258446 0 258502 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 260378 0 260434 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 262310 0 262366 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 1490 0 1546 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 320000 440000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 135500046
string GDS_FILE /home/htamas/progs/unigate-sky-comb/openlane/unigate/runs/22_12_11_19_17/results/signoff/unigate.magic.gds
string GDS_START 1678050
<< end >>

