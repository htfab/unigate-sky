module u31_ref (
    input [7:0] func,
    input [2:0] pin,
    output [2:0] wiring
);

reg [17:0] w;
assign wiring = w[3*pin+:3];

always @ (func) begin
    case (func)
        8'b00000000 : w = 18'b000_000_000_000_000_000;
        8'b00000001 : w = 18'b100_010_011_010_001_001;
        8'b00000010 : w = 18'b001_100_011_000_010_010;
        8'b00000011 : w = 18'b001_100_011_000_000_000;
        8'b00000100 : w = 18'b100_010_000_011_011_010;
        8'b00000101 : w = 18'b001_100_010_000_000_000;
        8'b00000110 : w = 18'b001_100_011_010_010_000;
        8'b00000111 : w = 18'b010_011_001_100_010_001;
        8'b00001000 : w = 18'b011_010_100_010_000_000;
        8'b00001001 : w = 18'b011_011_010_100_001_001;
        8'b00001010 : w = 18'b010_100_000_000_000_000;
        8'b00001011 : w = 18'b010_100_000_011_011_000;
        8'b00001100 : w = 18'b011_100_000_000_000_000;
        8'b00001101 : w = 18'b011_100_000_010_010_000;
        8'b00001110 : w = 18'b011_100_011_010_010_000;
        8'b00001111 : w = 18'b000_100_000_000_000_000;
        8'b00010000 : w = 18'b011_010_000_100_100_010;
        8'b00010001 : w = 18'b001_011_010_000_000_000;
        8'b00010010 : w = 18'b001_011_100_010_010_000;
        8'b00010011 : w = 18'b010_100_001_011_010_001;
        8'b00010100 : w = 18'b001_010_100_011_011_000;
        8'b00010101 : w = 18'b011_100_001_010_011_001;
        8'b00010110 : w = 18'b100_011_010_000_011_010;
        8'b00010111 : w = 18'b011_100_001_011_010_001;
        8'b00011000 : w = 18'b100_011_001_000_010_001;
        8'b00011001 : w = 18'b011_010_100_000_010_000;
        8'b00011010 : w = 18'b001_010_011_100_000_000;
        8'b00011011 : w = 18'b011_100_001_001_010_001;
        8'b00011100 : w = 18'b001_011_010_100_000_000;
        8'b00011101 : w = 18'b010_100_001_001_011_001;
        8'b00011110 : w = 18'b011_011_100_010_010_000;
        8'b00011111 : w = 18'b011_010_000_100_010_000;
        8'b00100000 : w = 18'b100_010_011_010_000_000;
        8'b00100001 : w = 18'b100_100_010_011_001_001;
        8'b00100010 : w = 18'b010_011_000_000_000_000;
        8'b00100011 : w = 18'b010_011_000_100_100_000;
        8'b00100100 : w = 18'b011_100_001_000_010_001;
        8'b00100101 : w = 18'b100_010_011_000_010_000;
        8'b00100110 : w = 18'b001_010_100_011_000_000;
        8'b00100111 : w = 18'b100_011_001_001_010_001;
        8'b00101000 : w = 18'b000_000_010_100_011_010;
        8'b00101001 : w = 18'b100_011_001_010_011_001;
        8'b00101010 : w = 18'b010_100_011_011_011_000;
        8'b00101011 : w = 18'b010_100_011_000_000_000;
        8'b00101100 : w = 18'b010_011_000_100_000_000;
        8'b00101101 : w = 18'b010_011_000_000_100_000;
        8'b00101110 : w = 18'b010_010_100_011_000_000;
        8'b00101111 : w = 18'b010_000_011_100_000_000;
        8'b00110000 : w = 18'b100_011_000_000_000_000;
        8'b00110001 : w = 18'b100_011_000_010_010_000;
        8'b00110010 : w = 18'b100_011_011_010_010_000;
        8'b00110011 : w = 18'b000_011_000_000_000_000;
        8'b00110100 : w = 18'b001_100_010_011_000_000;
        8'b00110101 : w = 18'b010_011_001_001_100_001;
        8'b00110110 : w = 18'b100_100_011_010_010_000;
        8'b00110111 : w = 18'b100_010_000_011_010_000;
        8'b00111000 : w = 18'b010_100_000_011_000_000;
        8'b00111001 : w = 18'b010_100_000_000_011_000;
        8'b00111010 : w = 18'b010_010_011_100_000_000;
        8'b00111011 : w = 18'b010_000_100_011_000_000;
        8'b00111100 : w = 18'b000_100_000_011_000_000;
        8'b00111101 : w = 18'b010_100_010_000_011_000;
        8'b00111110 : w = 18'b100_001_010_011_001_000;
        8'b00111111 : w = 18'b000_100_011_000_000_000;
        8'b01000000 : w = 18'b100_011_010_011_000_000;
        8'b01000001 : w = 18'b100_100_011_010_001_001;
        8'b01000010 : w = 18'b010_100_001_000_011_001;
        8'b01000011 : w = 18'b100_011_010_000_011_000;
        8'b01000100 : w = 18'b011_010_000_000_000_000;
        8'b01000101 : w = 18'b011_010_000_100_100_000;
        8'b01000110 : w = 18'b001_011_100_010_000_000;
        8'b01000111 : w = 18'b100_010_001_001_011_001;
        8'b01001000 : w = 18'b000_000_011_100_010_011;
        8'b01001001 : w = 18'b100_010_001_011_010_001;
        8'b01001010 : w = 18'b011_010_000_100_000_000;
        8'b01001011 : w = 18'b011_010_000_000_100_000;
        8'b01001100 : w = 18'b011_100_010_010_010_000;
        8'b01001101 : w = 18'b011_100_010_000_000_000;
        8'b01001110 : w = 18'b011_011_100_010_000_000;
        8'b01001111 : w = 18'b011_000_010_100_000_000;
        8'b01010000 : w = 18'b100_010_000_000_000_000;
        8'b01010001 : w = 18'b100_010_000_011_011_000;
        8'b01010010 : w = 18'b001_100_011_010_000_000;
        8'b01010011 : w = 18'b011_010_001_001_100_001;
        8'b01010100 : w = 18'b100_001_011_001_010_000;
        8'b01010101 : w = 18'b000_010_000_000_000_000;
        8'b01010110 : w = 18'b100_011_010_010_011_000;
        8'b01010111 : w = 18'b001_100_011_000_010_000;
        8'b01011000 : w = 18'b011_100_000_010_000_000;
        8'b01011001 : w = 18'b011_100_000_000_010_000;
        8'b01011010 : w = 18'b000_100_000_010_000_000;
        8'b01011011 : w = 18'b011_100_011_000_010_000;
        8'b01011100 : w = 18'b011_011_010_100_000_000;
        8'b01011101 : w = 18'b011_000_100_010_000_000;
        8'b01011110 : w = 18'b100_001_011_010_001_000;
        8'b01011111 : w = 18'b000_100_010_000_000_000;
        8'b01100000 : w = 18'b000_000_100_011_010_100;
        8'b01100001 : w = 18'b011_010_001_100_010_001;
        8'b01100010 : w = 18'b100_010_000_011_000_000;
        8'b01100011 : w = 18'b100_010_000_000_011_000;
        8'b01100100 : w = 18'b100_011_000_010_000_000;
        8'b01100101 : w = 18'b100_011_000_000_010_000;
        8'b01100110 : w = 18'b000_011_000_010_000_000;
        8'b01100111 : w = 18'b100_011_011_000_010_000;
        8'b01101000 : w = 18'b011_100_010_011_010_000;
        8'b01101001 : w = 18'b000_100_000_011_010_000;
        8'b01101010 : w = 18'b001_100_001_010_011_000;
        8'b01101011 : w = 18'b011_100_000_010_011_000;
        8'b01101100 : w = 18'b001_100_001_011_010_000;
        8'b01101101 : w = 18'b010_100_000_011_010_000;
        8'b01101110 : w = 18'b000_011_100_010_000_000;
        8'b01101111 : w = 18'b000_000_100_011_010_000;
        8'b01110000 : w = 18'b100_011_010_010_010_000;
        8'b01110001 : w = 18'b100_011_010_000_000_000;
        8'b01110010 : w = 18'b100_100_011_010_000_000;
        8'b01110011 : w = 18'b100_000_010_011_000_000;
        8'b01110100 : w = 18'b100_100_010_011_000_000;
        8'b01110101 : w = 18'b100_000_011_010_000_000;
        8'b01110110 : w = 18'b011_001_100_010_001_000;
        8'b01110111 : w = 18'b000_011_010_000_000_000;
        8'b01111000 : w = 18'b001_011_001_100_010_000;
        8'b01111001 : w = 18'b000_100_010_011_010_000;
        8'b01111010 : w = 18'b000_100_011_010_000_000;
        8'b01111011 : w = 18'b000_000_011_100_010_000;
        8'b01111100 : w = 18'b000_100_010_011_000_000;
        8'b01111101 : w = 18'b000_000_010_100_011_000;
        8'b01111110 : w = 18'b010_010_100_011_010_000;
        8'b01111111 : w = 18'b010_100_011_000_010_000;
        8'b10000000 : w = 18'b010_100_011_000_010_001;
        8'b10000001 : w = 18'b010_010_100_011_010_001;
        8'b10000010 : w = 18'b000_000_010_100_011_001;
        8'b10000011 : w = 18'b000_100_010_011_000_001;
        8'b10000100 : w = 18'b000_000_011_100_010_001;
        8'b10000101 : w = 18'b000_100_011_010_000_001;
        8'b10000110 : w = 18'b011_001_010_010_100_000;
        8'b10000111 : w = 18'b011_001_000_010_100_000;
        8'b10001000 : w = 18'b011_001_000_010_000_000;
        8'b10001001 : w = 18'b011_001_100_010_001_001;
        8'b10001010 : w = 18'b011_001_100_010_000_000;
        8'b10001011 : w = 18'b100_100_010_011_000_001;
        8'b10001100 : w = 18'b010_001_100_011_000_000;
        8'b10001101 : w = 18'b100_100_011_010_000_001;
        8'b10001110 : w = 18'b011_010_001_010_100_000;
        8'b10001111 : w = 18'b100_011_010_010_010_001;
        8'b10010000 : w = 18'b000_000_100_011_010_001;
        8'b10010001 : w = 18'b000_011_100_010_000_001;
        8'b10010010 : w = 18'b100_001_010_010_011_000;
        8'b10010011 : w = 18'b100_001_000_010_011_000;
        8'b10010100 : w = 18'b100_001_010_011_010_000;
        8'b10010101 : w = 18'b100_001_000_011_010_000;
        8'b10010110 : w = 18'b000_100_000_011_010_001;
        8'b10010111 : w = 18'b011_100_010_011_010_001;
        8'b10011000 : w = 18'b010_011_100_010_001_000;
        8'b10011001 : w = 18'b000_011_000_010_001_000;
        8'b10011010 : w = 18'b100_011_011_010_001_000;
        8'b10011011 : w = 18'b100_011_000_010_001_000;
        8'b10011100 : w = 18'b100_010_010_011_001_000;
        8'b10011101 : w = 18'b000_011_100_010_001_000;
        8'b10011110 : w = 18'b011_010_001_100_010_000;
        8'b10011111 : w = 18'b010_011_001_001_100_010;
        8'b10100000 : w = 18'b100_001_000_010_000_000;
        8'b10100001 : w = 18'b100_001_011_010_001_001;
        8'b10100010 : w = 18'b100_001_011_010_000_000;
        8'b10100011 : w = 18'b011_011_010_100_000_001;
        8'b10100100 : w = 18'b010_100_011_010_001_000;
        8'b10100101 : w = 18'b000_100_000_010_001_000;
        8'b10100110 : w = 18'b011_100_011_010_001_000;
        8'b10100111 : w = 18'b011_100_000_010_001_000;
        8'b10101000 : w = 18'b001_100_011_000_010_001;
        8'b10101001 : w = 18'b100_011_010_010_011_001;
        8'b10101010 : w = 18'b010_001_000_000_000_000;
        8'b10101011 : w = 18'b100_001_011_001_010_001;
        8'b10101100 : w = 18'b011_010_001_001_100_000;
        8'b10101101 : w = 18'b001_100_011_010_000_001;
        8'b10101110 : w = 18'b001_100_011_010_001_000;
        8'b10101111 : w = 18'b010_100_001_000_000_000;
        8'b10110000 : w = 18'b010_001_011_100_000_000;
        8'b10110001 : w = 18'b011_011_100_010_000_001;
        8'b10110010 : w = 18'b100_010_001_010_011_000;
        8'b10110011 : w = 18'b011_100_010_010_010_001;
        8'b10110100 : w = 18'b011_010_010_100_001_000;
        8'b10110101 : w = 18'b000_100_011_010_001_000;
        8'b10110110 : w = 18'b100_010_001_011_010_000;
        8'b10110111 : w = 18'b010_100_001_001_011_010;
        8'b10111000 : w = 18'b100_010_001_001_011_000;
        8'b10111001 : w = 18'b001_011_100_010_000_001;
        8'b10111010 : w = 18'b100_000_011_010_001_000;
        8'b10111011 : w = 18'b010_011_001_000_000_000;
        8'b10111100 : w = 18'b010_100_001_011_000_000;
        8'b10111101 : w = 18'b010_100_001_000_011_000;
        8'b10111110 : w = 18'b100_100_011_010_001_000;
        8'b10111111 : w = 18'b100_011_010_011_000_001;
        8'b11000000 : w = 18'b100_001_000_011_000_000;
        8'b11000001 : w = 18'b100_001_010_011_001_001;
        8'b11000010 : w = 18'b011_100_010_011_001_000;
        8'b11000011 : w = 18'b000_100_000_011_001_000;
        8'b11000100 : w = 18'b100_001_010_011_000_000;
        8'b11000101 : w = 18'b010_010_011_100_000_001;
        8'b11000110 : w = 18'b010_100_010_011_001_000;
        8'b11000111 : w = 18'b010_100_000_011_001_000;
        8'b11001000 : w = 18'b100_010_000_011_010_001;
        8'b11001001 : w = 18'b100_100_011_010_010_001;
        8'b11001010 : w = 18'b010_011_001_001_100_000;
        8'b11001011 : w = 18'b001_100_010_011_000_001;
        8'b11001100 : w = 18'b011_001_000_000_000_000;
        8'b11001101 : w = 18'b100_011_011_010_010_001;
        8'b11001110 : w = 18'b001_100_010_011_001_000;
        8'b11001111 : w = 18'b011_100_001_000_000_000;
        8'b11010000 : w = 18'b011_001_010_100_000_000;
        8'b11010001 : w = 18'b010_010_100_011_000_001;
        8'b11010010 : w = 18'b010_011_010_100_001_000;
        8'b11010011 : w = 18'b000_100_010_011_001_000;
        8'b11010100 : w = 18'b100_011_001_011_010_000;
        8'b11010101 : w = 18'b010_100_011_011_011_001;
        8'b11010110 : w = 18'b100_011_001_010_011_000;
        8'b11010111 : w = 18'b011_100_001_001_010_011;
        8'b11011000 : w = 18'b100_011_001_001_010_000;
        8'b11011001 : w = 18'b001_010_100_011_000_001;
        8'b11011010 : w = 18'b011_100_001_010_000_000;
        8'b11011011 : w = 18'b011_100_001_000_010_000;
        8'b11011100 : w = 18'b100_000_010_011_001_000;
        8'b11011101 : w = 18'b011_010_001_000_000_000;
        8'b11011110 : w = 18'b100_100_010_011_001_000;
        8'b11011111 : w = 18'b100_010_011_010_000_001;
        8'b11100000 : w = 18'b011_010_000_100_010_001;
        8'b11100001 : w = 18'b011_011_100_010_010_001;
        8'b11100010 : w = 18'b010_100_001_001_011_000;
        8'b11100011 : w = 18'b001_011_010_100_000_001;
        8'b11100100 : w = 18'b011_100_001_001_010_000;
        8'b11100101 : w = 18'b001_010_011_100_000_001;
        8'b11100110 : w = 18'b100_011_001_010_000_000;
        8'b11100111 : w = 18'b100_011_001_000_010_000;
        8'b11101000 : w = 18'b011_100_001_011_010_000;
        8'b11101001 : w = 18'b010_100_001_011_000_010;
        8'b11101010 : w = 18'b011_100_001_010_011_000;
        8'b11101011 : w = 18'b000_010_001_100_011_000;
        8'b11101100 : w = 18'b010_100_001_011_010_000;
        8'b11101101 : w = 18'b000_011_001_100_010_000;
        8'b11101110 : w = 18'b000_011_001_010_000_000;
        8'b11101111 : w = 18'b100_000_011_010_001_010;
        8'b11110000 : w = 18'b100_001_000_000_000_000;
        8'b11110001 : w = 18'b011_100_011_010_010_001;
        8'b11110010 : w = 18'b001_011_010_100_001_000;
        8'b11110011 : w = 18'b100_011_001_000_000_000;
        8'b11110100 : w = 18'b011_000_010_100_001_000;
        8'b11110101 : w = 18'b100_010_001_000_000_000;
        8'b11110110 : w = 18'b011_011_010_100_001_000;
        8'b11110111 : w = 18'b011_010_100_010_000_001;
        8'b11111000 : w = 18'b010_011_001_100_010_000;
        8'b11111001 : w = 18'b000_100_001_011_010_000;
        8'b11111010 : w = 18'b000_100_001_010_000_000;
        8'b11111011 : w = 18'b001_100_011_010_001_010;
        8'b11111100 : w = 18'b000_100_001_011_000_000;
        8'b11111101 : w = 18'b001_100_010_011_001_011;
        8'b11111110 : w = 18'b100_010_011_010_001_000;
        8'b11111111 : w = 18'b000_001_000_000_000_000;
    endcase
end

endmodule

