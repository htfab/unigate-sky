module u31_ref_tb ();

integer i;
reg [23:0] func;
wire [2:0] pin = i;
reg [17:0] wiring;
wire [2:0] wtest;
wire [7:0] fcmp = {func[21], func[18], func[15], func[12], func[9], func[6], func[3], func[0]};
wire [15:0] fres = {func[23], func[22], func[20], func[19], func[17], func[16], func[14], func[13],
                    func[11], func[10], func[8], func[7], func[5], func[4], func[2], func[1]};
wire assert = (wiring[3*i+:3] == wtest) && (fres == 16'b0);

wire [2:0] O = 3'b000;
wire [2:0] I = 3'b001;
wire [2:0] a = 3'b010;
wire [2:0] b = 3'b011;
wire [2:0] c = 3'b100;

u31_ref dut (
    .func(fcmp),
    .pin(pin),
    .wiring(wtest)
);

initial begin
    for (i=0; i<6; i=i+1) begin
        #1 func = {O, O, O, O, O, O, O, O}; wiring = {O, O, O, O, O, O}; #1 $display(assert);
        #1 func = {O, O, O, O, O, O, O, I}; wiring = {c, a, b, a, I, I}; #1 $display(assert);
        #1 func = {O, O, O, O, O, O, I, O}; wiring = {I, c, b, O, a, a}; #1 $display(assert);
        #1 func = {O, O, O, O, O, O, I, I}; wiring = {I, c, b, O, O, O}; #1 $display(assert);
        #1 func = {O, O, O, O, O, I, O, O}; wiring = {c, a, O, b, b, a}; #1 $display(assert);
        #1 func = {O, O, O, O, O, I, O, I}; wiring = {I, c, a, O, O, O}; #1 $display(assert);
        #1 func = {O, O, O, O, O, I, I, O}; wiring = {I, c, b, a, a, O}; #1 $display(assert);
        #1 func = {O, O, O, O, O, I, I, I}; wiring = {a, b, I, c, a, I}; #1 $display(assert);
        #1 func = {O, O, O, O, I, O, O, O}; wiring = {b, a, c, a, O, O}; #1 $display(assert);
        #1 func = {O, O, O, O, I, O, O, I}; wiring = {b, b, a, c, I, I}; #1 $display(assert);
        #1 func = {O, O, O, O, I, O, I, O}; wiring = {a, c, O, O, O, O}; #1 $display(assert);
        #1 func = {O, O, O, O, I, O, I, I}; wiring = {a, c, O, b, b, O}; #1 $display(assert);
        #1 func = {O, O, O, O, I, I, O, O}; wiring = {b, c, O, O, O, O}; #1 $display(assert);
        #1 func = {O, O, O, O, I, I, O, I}; wiring = {b, c, O, a, a, O}; #1 $display(assert);
        #1 func = {O, O, O, O, I, I, I, O}; wiring = {b, c, b, a, a, O}; #1 $display(assert);
        #1 func = {O, O, O, O, I, I, I, I}; wiring = {O, c, O, O, O, O}; #1 $display(assert);
        #1 func = {O, O, O, I, O, O, O, O}; wiring = {b, a, O, c, c, a}; #1 $display(assert);
        #1 func = {O, O, O, I, O, O, O, I}; wiring = {I, b, a, O, O, O}; #1 $display(assert);
        #1 func = {O, O, O, I, O, O, I, O}; wiring = {I, b, c, a, a, O}; #1 $display(assert);
        #1 func = {O, O, O, I, O, O, I, I}; wiring = {a, c, I, b, a, I}; #1 $display(assert);
        #1 func = {O, O, O, I, O, I, O, O}; wiring = {I, a, c, b, b, O}; #1 $display(assert);
        #1 func = {O, O, O, I, O, I, O, I}; wiring = {b, c, I, a, b, I}; #1 $display(assert);
        #1 func = {O, O, O, I, O, I, I, O}; wiring = {c, b, a, O, b, a}; #1 $display(assert);
        #1 func = {O, O, O, I, O, I, I, I}; wiring = {b, c, I, b, a, I}; #1 $display(assert);
        #1 func = {O, O, O, I, I, O, O, O}; wiring = {c, b, I, O, a, I}; #1 $display(assert);
        #1 func = {O, O, O, I, I, O, O, I}; wiring = {b, a, c, O, a, O}; #1 $display(assert);
        #1 func = {O, O, O, I, I, O, I, O}; wiring = {I, a, b, c, O, O}; #1 $display(assert);
        #1 func = {O, O, O, I, I, O, I, I}; wiring = {b, c, I, I, a, I}; #1 $display(assert);
        #1 func = {O, O, O, I, I, I, O, O}; wiring = {I, b, a, c, O, O}; #1 $display(assert);
        #1 func = {O, O, O, I, I, I, O, I}; wiring = {a, c, I, I, b, I}; #1 $display(assert);
        #1 func = {O, O, O, I, I, I, I, O}; wiring = {b, b, c, a, a, O}; #1 $display(assert);
        #1 func = {O, O, O, I, I, I, I, I}; wiring = {b, a, O, c, a, O}; #1 $display(assert);
        #1 func = {O, O, I, O, O, O, O, O}; wiring = {c, a, b, a, O, O}; #1 $display(assert);
        #1 func = {O, O, I, O, O, O, O, I}; wiring = {c, c, a, b, I, I}; #1 $display(assert);
        #1 func = {O, O, I, O, O, O, I, O}; wiring = {a, b, O, O, O, O}; #1 $display(assert);
        #1 func = {O, O, I, O, O, O, I, I}; wiring = {a, b, O, c, c, O}; #1 $display(assert);
        #1 func = {O, O, I, O, O, I, O, O}; wiring = {b, c, I, O, a, I}; #1 $display(assert);
        #1 func = {O, O, I, O, O, I, O, I}; wiring = {c, a, b, O, a, O}; #1 $display(assert);
        #1 func = {O, O, I, O, O, I, I, O}; wiring = {I, a, c, b, O, O}; #1 $display(assert);
        #1 func = {O, O, I, O, O, I, I, I}; wiring = {c, b, I, I, a, I}; #1 $display(assert);
        #1 func = {O, O, I, O, I, O, O, O}; wiring = {O, O, a, c, b, a}; #1 $display(assert);
        #1 func = {O, O, I, O, I, O, O, I}; wiring = {c, b, I, a, b, I}; #1 $display(assert);
        #1 func = {O, O, I, O, I, O, I, O}; wiring = {a, c, b, b, b, O}; #1 $display(assert);
        #1 func = {O, O, I, O, I, O, I, I}; wiring = {a, c, b, O, O, O}; #1 $display(assert);
        #1 func = {O, O, I, O, I, I, O, O}; wiring = {a, b, O, c, O, O}; #1 $display(assert);
        #1 func = {O, O, I, O, I, I, O, I}; wiring = {a, b, O, O, c, O}; #1 $display(assert);
        #1 func = {O, O, I, O, I, I, I, O}; wiring = {a, a, c, b, O, O}; #1 $display(assert);
        #1 func = {O, O, I, O, I, I, I, I}; wiring = {a, O, b, c, O, O}; #1 $display(assert);
        #1 func = {O, O, I, I, O, O, O, O}; wiring = {c, b, O, O, O, O}; #1 $display(assert);
        #1 func = {O, O, I, I, O, O, O, I}; wiring = {c, b, O, a, a, O}; #1 $display(assert);
        #1 func = {O, O, I, I, O, O, I, O}; wiring = {c, b, b, a, a, O}; #1 $display(assert);
        #1 func = {O, O, I, I, O, O, I, I}; wiring = {O, b, O, O, O, O}; #1 $display(assert);
        #1 func = {O, O, I, I, O, I, O, O}; wiring = {I, c, a, b, O, O}; #1 $display(assert);
        #1 func = {O, O, I, I, O, I, O, I}; wiring = {a, b, I, I, c, I}; #1 $display(assert);
        #1 func = {O, O, I, I, O, I, I, O}; wiring = {c, c, b, a, a, O}; #1 $display(assert);
        #1 func = {O, O, I, I, O, I, I, I}; wiring = {c, a, O, b, a, O}; #1 $display(assert);
        #1 func = {O, O, I, I, I, O, O, O}; wiring = {a, c, O, b, O, O}; #1 $display(assert);
        #1 func = {O, O, I, I, I, O, O, I}; wiring = {a, c, O, O, b, O}; #1 $display(assert);
        #1 func = {O, O, I, I, I, O, I, O}; wiring = {a, a, b, c, O, O}; #1 $display(assert);
        #1 func = {O, O, I, I, I, O, I, I}; wiring = {a, O, c, b, O, O}; #1 $display(assert);
        #1 func = {O, O, I, I, I, I, O, O}; wiring = {O, c, O, b, O, O}; #1 $display(assert);
        #1 func = {O, O, I, I, I, I, O, I}; wiring = {a, c, a, O, b, O}; #1 $display(assert);
        #1 func = {O, O, I, I, I, I, I, O}; wiring = {c, I, a, b, I, O}; #1 $display(assert);
        #1 func = {O, O, I, I, I, I, I, I}; wiring = {O, c, b, O, O, O}; #1 $display(assert);
        #1 func = {O, I, O, O, O, O, O, O}; wiring = {c, b, a, b, O, O}; #1 $display(assert);
        #1 func = {O, I, O, O, O, O, O, I}; wiring = {c, c, b, a, I, I}; #1 $display(assert);
        #1 func = {O, I, O, O, O, O, I, O}; wiring = {a, c, I, O, b, I}; #1 $display(assert);
        #1 func = {O, I, O, O, O, O, I, I}; wiring = {c, b, a, O, b, O}; #1 $display(assert);
        #1 func = {O, I, O, O, O, I, O, O}; wiring = {b, a, O, O, O, O}; #1 $display(assert);
        #1 func = {O, I, O, O, O, I, O, I}; wiring = {b, a, O, c, c, O}; #1 $display(assert);
        #1 func = {O, I, O, O, O, I, I, O}; wiring = {I, b, c, a, O, O}; #1 $display(assert);
        #1 func = {O, I, O, O, O, I, I, I}; wiring = {c, a, I, I, b, I}; #1 $display(assert);
        #1 func = {O, I, O, O, I, O, O, O}; wiring = {O, O, b, c, a, b}; #1 $display(assert);
        #1 func = {O, I, O, O, I, O, O, I}; wiring = {c, a, I, b, a, I}; #1 $display(assert);
        #1 func = {O, I, O, O, I, O, I, O}; wiring = {b, a, O, c, O, O}; #1 $display(assert);
        #1 func = {O, I, O, O, I, O, I, I}; wiring = {b, a, O, O, c, O}; #1 $display(assert);
        #1 func = {O, I, O, O, I, I, O, O}; wiring = {b, c, a, a, a, O}; #1 $display(assert);
        #1 func = {O, I, O, O, I, I, O, I}; wiring = {b, c, a, O, O, O}; #1 $display(assert);
        #1 func = {O, I, O, O, I, I, I, O}; wiring = {b, b, c, a, O, O}; #1 $display(assert);
        #1 func = {O, I, O, O, I, I, I, I}; wiring = {b, O, a, c, O, O}; #1 $display(assert);
        #1 func = {O, I, O, I, O, O, O, O}; wiring = {c, a, O, O, O, O}; #1 $display(assert);
        #1 func = {O, I, O, I, O, O, O, I}; wiring = {c, a, O, b, b, O}; #1 $display(assert);
        #1 func = {O, I, O, I, O, O, I, O}; wiring = {I, c, b, a, O, O}; #1 $display(assert);
        #1 func = {O, I, O, I, O, O, I, I}; wiring = {b, a, I, I, c, I}; #1 $display(assert);
        #1 func = {O, I, O, I, O, I, O, O}; wiring = {c, I, b, I, a, O}; #1 $display(assert);
        #1 func = {O, I, O, I, O, I, O, I}; wiring = {O, a, O, O, O, O}; #1 $display(assert);
        #1 func = {O, I, O, I, O, I, I, O}; wiring = {c, b, a, a, b, O}; #1 $display(assert);
        #1 func = {O, I, O, I, O, I, I, I}; wiring = {I, c, b, O, a, O}; #1 $display(assert);
        #1 func = {O, I, O, I, I, O, O, O}; wiring = {b, c, O, a, O, O}; #1 $display(assert);
        #1 func = {O, I, O, I, I, O, O, I}; wiring = {b, c, O, O, a, O}; #1 $display(assert);
        #1 func = {O, I, O, I, I, O, I, O}; wiring = {O, c, O, a, O, O}; #1 $display(assert);
        #1 func = {O, I, O, I, I, O, I, I}; wiring = {b, c, b, O, a, O}; #1 $display(assert);
        #1 func = {O, I, O, I, I, I, O, O}; wiring = {b, b, a, c, O, O}; #1 $display(assert);
        #1 func = {O, I, O, I, I, I, O, I}; wiring = {b, O, c, a, O, O}; #1 $display(assert);
        #1 func = {O, I, O, I, I, I, I, O}; wiring = {c, I, b, a, I, O}; #1 $display(assert);
        #1 func = {O, I, O, I, I, I, I, I}; wiring = {O, c, a, O, O, O}; #1 $display(assert);
        #1 func = {O, I, I, O, O, O, O, O}; wiring = {O, O, c, b, a, c}; #1 $display(assert);
        #1 func = {O, I, I, O, O, O, O, I}; wiring = {b, a, I, c, a, I}; #1 $display(assert);
        #1 func = {O, I, I, O, O, O, I, O}; wiring = {c, a, O, b, O, O}; #1 $display(assert);
        #1 func = {O, I, I, O, O, O, I, I}; wiring = {c, a, O, O, b, O}; #1 $display(assert);
        #1 func = {O, I, I, O, O, I, O, O}; wiring = {c, b, O, a, O, O}; #1 $display(assert);
        #1 func = {O, I, I, O, O, I, O, I}; wiring = {c, b, O, O, a, O}; #1 $display(assert);
        #1 func = {O, I, I, O, O, I, I, O}; wiring = {O, b, O, a, O, O}; #1 $display(assert);
        #1 func = {O, I, I, O, O, I, I, I}; wiring = {c, b, b, O, a, O}; #1 $display(assert);
        #1 func = {O, I, I, O, I, O, O, O}; wiring = {b, c, a, b, a, O}; #1 $display(assert);
        #1 func = {O, I, I, O, I, O, O, I}; wiring = {O, c, O, b, a, O}; #1 $display(assert);
        #1 func = {O, I, I, O, I, O, I, O}; wiring = {I, c, I, a, b, O}; #1 $display(assert);
        #1 func = {O, I, I, O, I, O, I, I}; wiring = {b, c, O, a, b, O}; #1 $display(assert);
        #1 func = {O, I, I, O, I, I, O, O}; wiring = {I, c, I, b, a, O}; #1 $display(assert);
        #1 func = {O, I, I, O, I, I, O, I}; wiring = {a, c, O, b, a, O}; #1 $display(assert);
        #1 func = {O, I, I, O, I, I, I, O}; wiring = {O, b, c, a, O, O}; #1 $display(assert);
        #1 func = {O, I, I, O, I, I, I, I}; wiring = {O, O, c, b, a, O}; #1 $display(assert);
        #1 func = {O, I, I, I, O, O, O, O}; wiring = {c, b, a, a, a, O}; #1 $display(assert);
        #1 func = {O, I, I, I, O, O, O, I}; wiring = {c, b, a, O, O, O}; #1 $display(assert);
        #1 func = {O, I, I, I, O, O, I, O}; wiring = {c, c, b, a, O, O}; #1 $display(assert);
        #1 func = {O, I, I, I, O, O, I, I}; wiring = {c, O, a, b, O, O}; #1 $display(assert);
        #1 func = {O, I, I, I, O, I, O, O}; wiring = {c, c, a, b, O, O}; #1 $display(assert);
        #1 func = {O, I, I, I, O, I, O, I}; wiring = {c, O, b, a, O, O}; #1 $display(assert);
        #1 func = {O, I, I, I, O, I, I, O}; wiring = {b, I, c, a, I, O}; #1 $display(assert);
        #1 func = {O, I, I, I, O, I, I, I}; wiring = {O, b, a, O, O, O}; #1 $display(assert);
        #1 func = {O, I, I, I, I, O, O, O}; wiring = {I, b, I, c, a, O}; #1 $display(assert);
        #1 func = {O, I, I, I, I, O, O, I}; wiring = {O, c, a, b, a, O}; #1 $display(assert);
        #1 func = {O, I, I, I, I, O, I, O}; wiring = {O, c, b, a, O, O}; #1 $display(assert);
        #1 func = {O, I, I, I, I, O, I, I}; wiring = {O, O, b, c, a, O}; #1 $display(assert);
        #1 func = {O, I, I, I, I, I, O, O}; wiring = {O, c, a, b, O, O}; #1 $display(assert);
        #1 func = {O, I, I, I, I, I, O, I}; wiring = {O, O, a, c, b, O}; #1 $display(assert);
        #1 func = {O, I, I, I, I, I, I, O}; wiring = {a, a, c, b, a, O}; #1 $display(assert);
        #1 func = {O, I, I, I, I, I, I, I}; wiring = {a, c, b, O, a, O}; #1 $display(assert);
        #1 func = {I, O, O, O, O, O, O, O}; wiring = {a, c, b, O, a, I}; #1 $display(assert);
        #1 func = {I, O, O, O, O, O, O, I}; wiring = {a, a, c, b, a, I}; #1 $display(assert);
        #1 func = {I, O, O, O, O, O, I, O}; wiring = {O, O, a, c, b, I}; #1 $display(assert);
        #1 func = {I, O, O, O, O, O, I, I}; wiring = {O, c, a, b, O, I}; #1 $display(assert);
        #1 func = {I, O, O, O, O, I, O, O}; wiring = {O, O, b, c, a, I}; #1 $display(assert);
        #1 func = {I, O, O, O, O, I, O, I}; wiring = {O, c, b, a, O, I}; #1 $display(assert);
        #1 func = {I, O, O, O, O, I, I, O}; wiring = {b, I, a, a, c, O}; #1 $display(assert);
        #1 func = {I, O, O, O, O, I, I, I}; wiring = {b, I, O, a, c, O}; #1 $display(assert);
        #1 func = {I, O, O, O, I, O, O, O}; wiring = {b, I, O, a, O, O}; #1 $display(assert);
        #1 func = {I, O, O, O, I, O, O, I}; wiring = {b, I, c, a, I, I}; #1 $display(assert);
        #1 func = {I, O, O, O, I, O, I, O}; wiring = {b, I, c, a, O, O}; #1 $display(assert);
        #1 func = {I, O, O, O, I, O, I, I}; wiring = {c, c, a, b, O, I}; #1 $display(assert);
        #1 func = {I, O, O, O, I, I, O, O}; wiring = {a, I, c, b, O, O}; #1 $display(assert);
        #1 func = {I, O, O, O, I, I, O, I}; wiring = {c, c, b, a, O, I}; #1 $display(assert);
        #1 func = {I, O, O, O, I, I, I, O}; wiring = {b, a, I, a, c, O}; #1 $display(assert);
        #1 func = {I, O, O, O, I, I, I, I}; wiring = {c, b, a, a, a, I}; #1 $display(assert);
        #1 func = {I, O, O, I, O, O, O, O}; wiring = {O, O, c, b, a, I}; #1 $display(assert);
        #1 func = {I, O, O, I, O, O, O, I}; wiring = {O, b, c, a, O, I}; #1 $display(assert);
        #1 func = {I, O, O, I, O, O, I, O}; wiring = {c, I, a, a, b, O}; #1 $display(assert);
        #1 func = {I, O, O, I, O, O, I, I}; wiring = {c, I, O, a, b, O}; #1 $display(assert);
        #1 func = {I, O, O, I, O, I, O, O}; wiring = {c, I, a, b, a, O}; #1 $display(assert);
        #1 func = {I, O, O, I, O, I, O, I}; wiring = {c, I, O, b, a, O}; #1 $display(assert);
        #1 func = {I, O, O, I, O, I, I, O}; wiring = {O, c, O, b, a, I}; #1 $display(assert);
        #1 func = {I, O, O, I, O, I, I, I}; wiring = {b, c, a, b, a, I}; #1 $display(assert);
        #1 func = {I, O, O, I, I, O, O, O}; wiring = {a, b, c, a, I, O}; #1 $display(assert);
        #1 func = {I, O, O, I, I, O, O, I}; wiring = {O, b, O, a, I, O}; #1 $display(assert);
        #1 func = {I, O, O, I, I, O, I, O}; wiring = {c, b, b, a, I, O}; #1 $display(assert);
        #1 func = {I, O, O, I, I, O, I, I}; wiring = {c, b, O, a, I, O}; #1 $display(assert);
        #1 func = {I, O, O, I, I, I, O, O}; wiring = {c, a, a, b, I, O}; #1 $display(assert);
        #1 func = {I, O, O, I, I, I, O, I}; wiring = {O, b, c, a, I, O}; #1 $display(assert);
        #1 func = {I, O, O, I, I, I, I, O}; wiring = {b, a, I, c, a, O}; #1 $display(assert);
        #1 func = {I, O, O, I, I, I, I, I}; wiring = {a, b, I, I, c, a}; #1 $display(assert);
        #1 func = {I, O, I, O, O, O, O, O}; wiring = {c, I, O, a, O, O}; #1 $display(assert);
        #1 func = {I, O, I, O, O, O, O, I}; wiring = {c, I, b, a, I, I}; #1 $display(assert);
        #1 func = {I, O, I, O, O, O, I, O}; wiring = {c, I, b, a, O, O}; #1 $display(assert);
        #1 func = {I, O, I, O, O, O, I, I}; wiring = {b, b, a, c, O, I}; #1 $display(assert);
        #1 func = {I, O, I, O, O, I, O, O}; wiring = {a, c, b, a, I, O}; #1 $display(assert);
        #1 func = {I, O, I, O, O, I, O, I}; wiring = {O, c, O, a, I, O}; #1 $display(assert);
        #1 func = {I, O, I, O, O, I, I, O}; wiring = {b, c, b, a, I, O}; #1 $display(assert);
        #1 func = {I, O, I, O, O, I, I, I}; wiring = {b, c, O, a, I, O}; #1 $display(assert);
        #1 func = {I, O, I, O, I, O, O, O}; wiring = {I, c, b, O, a, I}; #1 $display(assert);
        #1 func = {I, O, I, O, I, O, O, I}; wiring = {c, b, a, a, b, I}; #1 $display(assert);
        #1 func = {I, O, I, O, I, O, I, O}; wiring = {a, I, O, O, O, O}; #1 $display(assert);
        #1 func = {I, O, I, O, I, O, I, I}; wiring = {c, I, b, I, a, I}; #1 $display(assert);
        #1 func = {I, O, I, O, I, I, O, O}; wiring = {b, a, I, I, c, O}; #1 $display(assert);
        #1 func = {I, O, I, O, I, I, O, I}; wiring = {I, c, b, a, O, I}; #1 $display(assert);
        #1 func = {I, O, I, O, I, I, I, O}; wiring = {I, c, b, a, I, O}; #1 $display(assert);
        #1 func = {I, O, I, O, I, I, I, I}; wiring = {a, c, I, O, O, O}; #1 $display(assert);
        #1 func = {I, O, I, I, O, O, O, O}; wiring = {a, I, b, c, O, O}; #1 $display(assert);
        #1 func = {I, O, I, I, O, O, O, I}; wiring = {b, b, c, a, O, I}; #1 $display(assert);
        #1 func = {I, O, I, I, O, O, I, O}; wiring = {c, a, I, a, b, O}; #1 $display(assert);
        #1 func = {I, O, I, I, O, O, I, I}; wiring = {b, c, a, a, a, I}; #1 $display(assert);
        #1 func = {I, O, I, I, O, I, O, O}; wiring = {b, a, a, c, I, O}; #1 $display(assert);
        #1 func = {I, O, I, I, O, I, O, I}; wiring = {O, c, b, a, I, O}; #1 $display(assert);
        #1 func = {I, O, I, I, O, I, I, O}; wiring = {c, a, I, b, a, O}; #1 $display(assert);
        #1 func = {I, O, I, I, O, I, I, I}; wiring = {a, c, I, I, b, a}; #1 $display(assert);
        #1 func = {I, O, I, I, I, O, O, O}; wiring = {c, a, I, I, b, O}; #1 $display(assert);
        #1 func = {I, O, I, I, I, O, O, I}; wiring = {I, b, c, a, O, I}; #1 $display(assert);
        #1 func = {I, O, I, I, I, O, I, O}; wiring = {c, O, b, a, I, O}; #1 $display(assert);
        #1 func = {I, O, I, I, I, O, I, I}; wiring = {a, b, I, O, O, O}; #1 $display(assert);
        #1 func = {I, O, I, I, I, I, O, O}; wiring = {a, c, I, b, O, O}; #1 $display(assert);
        #1 func = {I, O, I, I, I, I, O, I}; wiring = {a, c, I, O, b, O}; #1 $display(assert);
        #1 func = {I, O, I, I, I, I, I, O}; wiring = {c, c, b, a, I, O}; #1 $display(assert);
        #1 func = {I, O, I, I, I, I, I, I}; wiring = {c, b, a, b, O, I}; #1 $display(assert);
        #1 func = {I, I, O, O, O, O, O, O}; wiring = {c, I, O, b, O, O}; #1 $display(assert);
        #1 func = {I, I, O, O, O, O, O, I}; wiring = {c, I, a, b, I, I}; #1 $display(assert);
        #1 func = {I, I, O, O, O, O, I, O}; wiring = {b, c, a, b, I, O}; #1 $display(assert);
        #1 func = {I, I, O, O, O, O, I, I}; wiring = {O, c, O, b, I, O}; #1 $display(assert);
        #1 func = {I, I, O, O, O, I, O, O}; wiring = {c, I, a, b, O, O}; #1 $display(assert);
        #1 func = {I, I, O, O, O, I, O, I}; wiring = {a, a, b, c, O, I}; #1 $display(assert);
        #1 func = {I, I, O, O, O, I, I, O}; wiring = {a, c, a, b, I, O}; #1 $display(assert);
        #1 func = {I, I, O, O, O, I, I, I}; wiring = {a, c, O, b, I, O}; #1 $display(assert);
        #1 func = {I, I, O, O, I, O, O, O}; wiring = {c, a, O, b, a, I}; #1 $display(assert);
        #1 func = {I, I, O, O, I, O, O, I}; wiring = {c, c, b, a, a, I}; #1 $display(assert);
        #1 func = {I, I, O, O, I, O, I, O}; wiring = {a, b, I, I, c, O}; #1 $display(assert);
        #1 func = {I, I, O, O, I, O, I, I}; wiring = {I, c, a, b, O, I}; #1 $display(assert);
        #1 func = {I, I, O, O, I, I, O, O}; wiring = {b, I, O, O, O, O}; #1 $display(assert);
        #1 func = {I, I, O, O, I, I, O, I}; wiring = {c, b, b, a, a, I}; #1 $display(assert);
        #1 func = {I, I, O, O, I, I, I, O}; wiring = {I, c, a, b, I, O}; #1 $display(assert);
        #1 func = {I, I, O, O, I, I, I, I}; wiring = {b, c, I, O, O, O}; #1 $display(assert);
        #1 func = {I, I, O, I, O, O, O, O}; wiring = {b, I, a, c, O, O}; #1 $display(assert);
        #1 func = {I, I, O, I, O, O, O, I}; wiring = {a, a, c, b, O, I}; #1 $display(assert);
        #1 func = {I, I, O, I, O, O, I, O}; wiring = {a, b, a, c, I, O}; #1 $display(assert);
        #1 func = {I, I, O, I, O, O, I, I}; wiring = {O, c, a, b, I, O}; #1 $display(assert);
        #1 func = {I, I, O, I, O, I, O, O}; wiring = {c, b, I, b, a, O}; #1 $display(assert);
        #1 func = {I, I, O, I, O, I, O, I}; wiring = {a, c, b, b, b, I}; #1 $display(assert);
        #1 func = {I, I, O, I, O, I, I, O}; wiring = {c, b, I, a, b, O}; #1 $display(assert);
        #1 func = {I, I, O, I, O, I, I, I}; wiring = {b, c, I, I, a, b}; #1 $display(assert);
        #1 func = {I, I, O, I, I, O, O, O}; wiring = {c, b, I, I, a, O}; #1 $display(assert);
        #1 func = {I, I, O, I, I, O, O, I}; wiring = {I, a, c, b, O, I}; #1 $display(assert);
        #1 func = {I, I, O, I, I, O, I, O}; wiring = {b, c, I, a, O, O}; #1 $display(assert);
        #1 func = {I, I, O, I, I, O, I, I}; wiring = {b, c, I, O, a, O}; #1 $display(assert);
        #1 func = {I, I, O, I, I, I, O, O}; wiring = {c, O, a, b, I, O}; #1 $display(assert);
        #1 func = {I, I, O, I, I, I, O, I}; wiring = {b, a, I, O, O, O}; #1 $display(assert);
        #1 func = {I, I, O, I, I, I, I, O}; wiring = {c, c, a, b, I, O}; #1 $display(assert);
        #1 func = {I, I, O, I, I, I, I, I}; wiring = {c, a, b, a, O, I}; #1 $display(assert);
        #1 func = {I, I, I, O, O, O, O, O}; wiring = {b, a, O, c, a, I}; #1 $display(assert);
        #1 func = {I, I, I, O, O, O, O, I}; wiring = {b, b, c, a, a, I}; #1 $display(assert);
        #1 func = {I, I, I, O, O, O, I, O}; wiring = {a, c, I, I, b, O}; #1 $display(assert);
        #1 func = {I, I, I, O, O, O, I, I}; wiring = {I, b, a, c, O, I}; #1 $display(assert);
        #1 func = {I, I, I, O, O, I, O, O}; wiring = {b, c, I, I, a, O}; #1 $display(assert);
        #1 func = {I, I, I, O, O, I, O, I}; wiring = {I, a, b, c, O, I}; #1 $display(assert);
        #1 func = {I, I, I, O, O, I, I, O}; wiring = {c, b, I, a, O, O}; #1 $display(assert);
        #1 func = {I, I, I, O, O, I, I, I}; wiring = {c, b, I, O, a, O}; #1 $display(assert);
        #1 func = {I, I, I, O, I, O, O, O}; wiring = {b, c, I, b, a, O}; #1 $display(assert);
        #1 func = {I, I, I, O, I, O, O, I}; wiring = {a, c, I, b, O, a}; #1 $display(assert);
        #1 func = {I, I, I, O, I, O, I, O}; wiring = {b, c, I, a, b, O}; #1 $display(assert);
        #1 func = {I, I, I, O, I, O, I, I}; wiring = {O, a, I, c, b, O}; #1 $display(assert);
        #1 func = {I, I, I, O, I, I, O, O}; wiring = {a, c, I, b, a, O}; #1 $display(assert);
        #1 func = {I, I, I, O, I, I, O, I}; wiring = {O, b, I, c, a, O}; #1 $display(assert);
        #1 func = {I, I, I, O, I, I, I, O}; wiring = {O, b, I, a, O, O}; #1 $display(assert);
        #1 func = {I, I, I, O, I, I, I, I}; wiring = {c, O, b, a, I, a}; #1 $display(assert);
        #1 func = {I, I, I, I, O, O, O, O}; wiring = {c, I, O, O, O, O}; #1 $display(assert);
        #1 func = {I, I, I, I, O, O, O, I}; wiring = {b, c, b, a, a, I}; #1 $display(assert);
        #1 func = {I, I, I, I, O, O, I, O}; wiring = {I, b, a, c, I, O}; #1 $display(assert);
        #1 func = {I, I, I, I, O, O, I, I}; wiring = {c, b, I, O, O, O}; #1 $display(assert);
        #1 func = {I, I, I, I, O, I, O, O}; wiring = {b, O, a, c, I, O}; #1 $display(assert);
        #1 func = {I, I, I, I, O, I, O, I}; wiring = {c, a, I, O, O, O}; #1 $display(assert);
        #1 func = {I, I, I, I, O, I, I, O}; wiring = {b, b, a, c, I, O}; #1 $display(assert);
        #1 func = {I, I, I, I, O, I, I, I}; wiring = {b, a, c, a, O, I}; #1 $display(assert);
        #1 func = {I, I, I, I, I, O, O, O}; wiring = {a, b, I, c, a, O}; #1 $display(assert);
        #1 func = {I, I, I, I, I, O, O, I}; wiring = {O, c, I, b, a, O}; #1 $display(assert);
        #1 func = {I, I, I, I, I, O, I, O}; wiring = {O, c, I, a, O, O}; #1 $display(assert);
        #1 func = {I, I, I, I, I, O, I, I}; wiring = {I, c, b, a, I, a}; #1 $display(assert);
        #1 func = {I, I, I, I, I, I, O, O}; wiring = {O, c, I, b, O, O}; #1 $display(assert);
        #1 func = {I, I, I, I, I, I, O, I}; wiring = {I, c, a, b, I, b}; #1 $display(assert);
        #1 func = {I, I, I, I, I, I, I, O}; wiring = {c, a, b, a, I, O}; #1 $display(assert);
        #1 func = {I, I, I, I, I, I, I, I}; wiring = {O, I, O, O, O, O}; #1 $display(assert);
    end
end

endmodule

